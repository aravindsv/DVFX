`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:28:46 03/02/2016 
// Design Name: 
// Module Name:    sinTable 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module sinTable(
    input clk,
    output [7:0] sFast,
    output [7:0] sMid,
    output [7:0] sSlow
    );


endmodule
